---------------------------------------------------
--Vinicius Malaman Soares
--Iowa State University
--Sep, 2024
---------------------------------------------------
--Test bench for a generic N-bit 2:1 Multiplexer
---------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;
library std;
use std.textio.all;

entity tb_N_bit_mux2t1 is
	generic(gCLK_HPER	: time := 10 ns);
end tb_N_bit_mux2t1;

architecture mixed of tb_N_bit_mux2t1 is


component mux2t1_N is
	generic(N: integer := 16);
	port(i_S	: in std_logic;
	     i_D0,i_D1  : in std_logic_vector(N-1 downto 0);
	     o_O	: out std_logic_vector(N-1 downto 0));
end component;

signal CLK, reset	: std_logic := '0';

constant N : integer := 16; -- Constant to be used as the N for testing purpose

signal s_D0	:std_logic_vector(N-1 downto 0);
signal s_D1   : std_logic_vector(N-1 downto 0) ;
signal s_S  : std_logic :='0';
signal s_O   : std_logic_vector(N-1 downto 0);

begin

	DUT0: mux2t1_N
	port map(i_D0=>s_D0,i_D1=>s_D1,i_S=>s_S,o_O=>s_O);

--first process is to setup the CLK
P_CLK: process
begin
	CLK<='1';
	wait for gCLK_HPER;
	CLK<= '0';
	wait for gCLK_HPER;
end process;
--second set the reset
P_RST: process
begin 
	reset<='0';
	wait for gCLK_HPER/2;
	reset<='1';
	wait for gCLK_HPER*2;
	reset <= '0';
	wait;
end process;

P_TEST_CASES: process
begin
	wait for gCLK_HPER/2;-- wait so the change doesnt happen at the edge

	--000
	G_Test1_Loop: for i in 0 to N-1 loop --loop through N-1 times and assign the vectors with either high or low
	s_S<='0';
	s_D0(i)<= '0';
	s_D1(i)<='0';
	end loop;
	wait for gCLK_HPER*2;
	--100
	G_Test2_Loop: for i in 0 to N-1 loop
 	s_S<='1';
	s_D1(i)<='0';
	s_D0(i)<= '0';
	end loop;
	wait for gCLK_HPER*2;
	--001
	G_Test3_Loop: for i in 0 to N-1 loop
 	s_S<='0';
	s_D1(i)<='0';
	s_D0(i)<= '1';
	end loop;
	wait for gCLK_HPER*2;
	--110
	G_Test4_Loop: for i in 0 to N-1 loop
 	s_S<='1';
	s_D1(i)<='1';
	s_D0(i)<= '0';
	end loop;
	wait for gCLK_HPER*2;
	
	
	--Special Tests
 	s_S<='0';
	s_D1<=x"F82C";
	s_D0<= x"AB9C";
	wait for gCLK_HPER*2;

	s_S<='1';
	s_D1<=x"F82C";
	s_D0<= x"AB9C";
	wait for gCLK_HPER*2;

	s_S<='0';
	s_D1<=x"F822";
	s_D0<= x"AFF1";
	wait for gCLK_HPER*2;

end process;


end mixed;


